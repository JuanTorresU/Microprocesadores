--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   16:41:28 11/09/2017
-- Design Name:   
-- Module Name:   C:/Proyectos ISE/Proyecto2/sim_1.vhd
-- Project Name:  Proyecto2
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: Memoria
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY sim_mem IS
END sim_mem;
 
ARCHITECTURE behavior OF sim_mem IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT Memoria
    PORT(
         a : IN  std_logic_vector(13 downto 0);
         d : IN  std_logic_vector(23 downto 0);
         dpra : IN  std_logic_vector(13 downto 0);
         clk : IN  std_logic;
         we : IN  std_logic;
         spo : OUT  std_logic_vector(23 downto 0);
         dpo : OUT  std_logic_vector(23 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal a : std_logic_vector(13 downto 0) := (others => '0');
   signal d : std_logic_vector(23 downto 0) := (others => '0');
   signal dpra : std_logic_vector(13 downto 0) := (others => '0');
   signal clk : std_logic := '0';
   signal we : std_logic := '0';

 	--Outputs
   signal spo : std_logic_vector(23 downto 0);
   signal dpo : std_logic_vector(23 downto 0);

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: Memoria PORT MAP (
          a => a,
          d => d,
          dpra => dpra,
          clk => clk,
          we => we,
          spo => spo,
          dpo => dpo
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	

      wait for clk_period*10;

      -- insert stimulus here 

      wait;
   end process;

END;
