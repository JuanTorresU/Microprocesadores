
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

entity RANDOM_CIRCUIT is
  port(
  
  );

end RANDOM_CIRCUIT;

architecture Behavioral of RANDOM_CIRCUIT is

begin

process()



end Behavioral;

